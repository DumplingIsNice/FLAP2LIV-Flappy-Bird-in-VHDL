--	GRAPHICS_PKG
--
--	Authors:		Callum McDowell, Hao Lin
--	Date:			May 2021
--	Course:		CS305 Miniproject
--
--
--	Summary
--
--		GRAPHICS_PKG is the shared format for sending, storing, and
--		accessing font render requests.
--
--		Each request is a packet of the form:
--		[col, row, scale, address, r, g, b]
--
--		col and row:	denote the top left corner of the font render (where to begin).
--		scale:			denotes what the bitmap should be multiplied by (at 1, 8x8 -> 8x8)
--		address:			is the address in CHAR_ROM ROM memory of the font 8x8 bitmap
--		r,g,b:			the colour the font should be rendered in (overrides previous values)
--
--		As VHDL synthesis has limited array dimension support we split the packet into
--		1D arrays of equal size (queue length), and access the relevant data in parallel.
--
--		Various other constants and records for the TRACKER, GENERATOR, and GRAPHICS_OBJECTS
--		are also stored here.


LIBRARY	IEEE;
USE		IEEE.STD_LOGIC_1164.all;
USE 		IEEE.NUMERIC_STD.all;

PACKAGE graphics_pkg IS

	-- GAMEPLAY MECHANICS CONSTANTS --
CONSTANT	DIFFICULTY_THRESHOLD_1		: UNSIGNED(7 downto 0)	:= TO_UNSIGNED(7,8);
CONSTANT DIFFICULTY_THRESHOLD_2		: UNSIGNED(7 downto 0)	:= TO_UNSIGNED(15,8);
CONSTANT DIFFICULTY_THRESHOLD_3		: UNSIGNED(7 downto 0)	:= TO_UNSIGNED(95,8);


	-- FONT --
	-- Break up font packet [col, row, scale, address] into 1D arrays for synthesis
CONSTANT FONT_QUEUE_LENGTH	: INTEGER := 23;

TYPE font_cols			IS ARRAY (FONT_QUEUE_LENGTH downto 0) OF STD_LOGIC_VECTOR(9 downto 0);
TYPE font_rows			IS ARRAY (FONT_QUEUE_LENGTH downto 0) OF STD_LOGIC_VECTOR(9 downto 0);
TYPE font_scales		IS ARRAY (FONT_QUEUE_LENGTH downto 0) OF STD_LOGIC_VECTOR(5 downto 0);
TYPE font_addresses	IS ARRAY (FONT_QUEUE_LENGTH downto 0) OF STD_LOGIC_VECTOR(5 downto 0);

SUBTYPE font_colour_packet IS STD_LOGIC_VECTOR(3 downto 0);
TYPE font_colour		IS ARRAY (FONT_QUEUE_LENGTH downto 0) OF FONT_COLOUR_PACKET;


	-- OBJECT --
	-- Each object queue has packets [col_left, row_upper, col_right, row_lower, type, r, g, b]
	-- left,upper describes the point the vector rectangle begins.
	-- right,lower describes the point the vector rectangle ends.
CONSTANT OBJ_QUEUE_LENGTH : INTEGER := 23;
	
TYPE obj_cols			IS ARRAY (OBJ_QUEUE_LENGTH downto 0) OF STD_LOGIC_VECTOR(9 downto 0);
TYPE obj_rows			IS ARRAY (OBJ_QUEUE_LENGTH downto 0) OF STD_LOGIC_VECTOR(9 downto 0);

SUBTYPE obj_type_packet IS STD_LOGIC_VECTOR(3 downto 0);
TYPE obj_types			IS ARRAY (OBJ_QUEUE_LENGTH downto 0) OF OBJ_TYPE_PACKET;
TYPE obj_colours		IS ARRAY (OBJ_QUEUE_LENGTH downto 0) OF FONT_COLOUR_PACKET;

TYPE obj_queue_packet IS RECORD
	-- record is used for structured storage in generator memory
	col					: STD_LOGIC_VECTOR(9 downto 0);
	row					: STD_LOGIC_VECTOR(9 downto 0);
	obj_type				: OBJ_TYPE_PACKET;
	r						: FONT_COLOUR_PACKET;
	g						: FONT_COLOUR_PACKET;
	b						: FONT_COLOUR_PACKET;
END RECORD obj_queue_packet;




	-- OBJECT HELPERS --
	-- (3, 2) = top coordinate (col, row), (1, 0) = bot coordinate (col, row)
TYPE obj_pos 			IS ARRAY (3 downto 0) OF STD_LOGIC_VECTOR (9 downto 0);
TYPE obj_mem 			IS ARRAY(OBJ_QUEUE_LENGTH downto 0) OF OBJ_POS;

CONSTANT OBJ_POS_ALL_ZERO 	: obj_pos 								:= (others => "0000000000");
CONSTANT OBJ_COLS_ALL_ZERO : obj_cols 								:= (others => "0000000000");
CONSTANT TEN_BIT_ALL_ZERO 	: STD_LOGIC_VECTOR (9 downto 0) 	:= "0000000000";
CONSTANT OBJ_COLOUR_ZERO	: FONT_COLOUR_PACKET					:= "0000";

CONSTANT GAP_FACTOR 			: STD_LOGIC_VECTOR(6 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(10, 7));
CONSTANT BORDER_MARGIN 		: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(40, 10));
CONSTANT GAP_HEIGHT 			: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(192, 10));

CONSTANT SCREEN_TOP			: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(0, 10));
CONSTANT SCREEN_BOT			: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(479, 10));
CONSTANT SCREEN_LEFT			: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(0, 10));
CONSTANT SCREEN_RIGHT		: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(639, 10));

CONSTANT PIPE_WIDTH 			: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(40, 10));
CONSTANT DIS_BETWEEN_PIPE 	: INTEGER := 320;
CONSTANT HALF_DIS_BETWEEN_PIPE 	: INTEGER := 160;

CONSTANT PIPE_TYPE			: OBJ_TYPE_PACKET						:= "0000";
CONSTANT PIPE_COLOUR			: FONT_COLOUR_PACKET					:= "0000";

CONSTANT BIRD_POSITION		: INTEGER								:= 200;

-- Pickup Positions
-- CONSTANT PICKUP_TOP_COL		: STD_LOGIC_VECTOR(9 downto 0)			:= STD_LOGIC_VECTOR(TO_UNSIGNED(32, 10));
CONSTANT PICKUP_TOP_ROW		: STD_LOGIC_VECTOR(9 downto 0)			:= STD_LOGIC_VECTOR(TO_UNSIGNED(32, 10));
-- CONSTANT PICKUP_BOT_COL		: STD_LOGIC_VECTOR(9 downto 0)			:= STD_LOGIC_VECTOR(TO_UNSIGNED(32, 10));
CONSTANT PICKUP_BOT_ROW		: STD_LOGIC_VECTOR(9 downto 0)			:= STD_LOGIC_VECTOR(TO_UNSIGNED(416, 10));

-- Chance is N out of 10.
CONSTANT INVI_CHANCE		: STD_LOGIC_VECTOR(3 downto 0)			:= STD_LOGIC_VECTOR(TO_UNSIGNED(3, 4));
CONSTANT INVI_TYPE			: OBJ_TYPE_PACKET						:= STD_LOGIC_VECTOR(TO_UNSIGNED(1, 4));
CONSTANT LIFE_CHANCE		: STD_LOGIC_VECTOR(3 downto 0)			:= STD_LOGIC_VECTOR(TO_UNSIGNED(3, 4));
CONSTANT LIFE_TYPE			: OBJ_TYPE_PACKET						:= STD_LOGIC_VECTOR(TO_UNSIGNED(2, 4));
CONSTANT COLOUR_SH_CHANCE	: STD_LOGIC_VECTOR(3 downto 0)			:= STD_LOGIC_VECTOR(TO_UNSIGNED(4, 4));
CONSTANT COLOUR_SH_TYPE		: OBJ_TYPE_PACKET						:= STD_LOGIC_VECTOR(TO_UNSIGNED(3, 4));

CONSTANT NULL_TYPE			: OBJ_TYPE_PACKET						:= "0000";

TYPE IS_SCORED_ARRAY		IS ARRAY (OBJ_QUEUE_LENGTH downto 0) OF STD_LOGIC;

CONSTANT DIFF_0 				: STD_LOGIC_VECTOR(1 downto 0)	:= "00";
CONSTANT DIFF_1 				: STD_LOGIC_VECTOR(1 downto 0)	:= "01";
CONSTANT DIFF_2 				: STD_LOGIC_VECTOR(1 downto 0)	:= "10";
CONSTANT DIFF_3 				: STD_LOGIC_VECTOR(1 downto 0)	:= "11";

CONSTANT DEFAULT_SPEED		: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(2, 10));
CONSTANT SPEED_1				: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(4, 10));
CONSTANT SPEED_2				: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(8, 10));
CONSTANT SPEED_3				: STD_LOGIC_VECTOR(9 downto 0)	:= STD_LOGIC_VECTOR(TO_UNSIGNED(16, 10));

CONSTANT UPPER_COLLISION	: UNSIGNED(9 downto 0)				:= TO_UNSIGNED(33,10);	-- 1/2 sprite height (i.e. 0.5*8*6) + 10px margin
CONSTANT LOWER_COLLISION	: UNSIGNED(9 downto 0)				:= TO_UNSIGNED(427,10);	-- 479 - sprite heigh (8*6) + 4px margin

	-- CONSTANTS --
CONSTANT CURSOR_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"77";
CONSTANT BIRD_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"76";

CONSTANT HEART_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"74";

CONSTANT A_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"01";
CONSTANT B_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"02";
CONSTANT C_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"03";
CONSTANT D_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"04";
CONSTANT E_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"05";
CONSTANT F_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"06";
CONSTANT G_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"07";
CONSTANT H_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"10";
CONSTANT I_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"11";
CONSTANT J_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"12";
CONSTANT K_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"13";
CONSTANT L_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"14";
CONSTANT M_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"15";
CONSTANT N_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"16";
CONSTANT O_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"17";
CONSTANT P_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"20";
CONSTANT Q_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"21";
CONSTANT R_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"22";
CONSTANT S_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"23";
CONSTANT T_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"24";
CONSTANT U_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"25";
CONSTANT V_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"26";
CONSTANT W_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"27";
CONSTANT X_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"30";
CONSTANT Y_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"31";
CONSTANT Z_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"32";
CONSTANT SPACE_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"40";

CONSTANT SQUARE_BRACKET_OPEN_ADDRESS	: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"33";
CONSTANT SQUARE_BRACKET_CLOSE_ADDRESS	: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"35";
CONSTANT DOWN_ARROW_ADDRESS				: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"34";
CONSTANT UP_ARROW_ADDRESS					: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"36";
CONSTANT RIGHT_ARROW_ADDRESS				: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"37";
CONSTANT ASTERISK_ADDRESS					: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"52";

CONSTANT ZERO_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"60";
CONSTANT ONE_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"61";
CONSTANT TWO_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"62";
CONSTANT THREE_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"63";
CONSTANT FOUR_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"64";
CONSTANT FIVE_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"65";
CONSTANT SIX_ADDRESS			: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"66";
CONSTANT SEVEN_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"67";
CONSTANT EIGHT_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"70";
CONSTANT NINE_ADDRESS		: STD_LOGIC_VECTOR (5 DOWNTO 0) := o"71";

END PACKAGE graphics_pkg;