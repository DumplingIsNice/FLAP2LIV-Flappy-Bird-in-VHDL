-- MAIN

-- Opening state machine for selecting a mode and beginning
-- Instigates gameplay loop.
